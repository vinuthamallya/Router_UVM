

typedef enum {BAD_XTN, GOOD_XTN}xtn_type;
